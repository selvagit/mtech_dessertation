// test project for revising the verilog

module  epcri_rx ( tx_payload_len, info_to_tx, data_to_mem, send_write_resp, sen_read_resp,
                    inp_clk, rx_buff, read_flg, reset);
input wire reset;
input wire[7:0] rx_buff;
input wire inp_clk;
input wire read_flg;
output wire send_write_resp;
output wire read_write_resp;
output reg[7:0] info_to_tx;

reg [7:0] inp_addr;
integer payload_len;

always @(posedge reset)
begin
    inp_addr <= 0;
    payload_len <= 0;
    send_write_resp <= 0;
    read_write_resp <= 0;
end

always @(posedge inp_clk)
begin
    if (read_flg)
    begin
        info_to_rx <= inp_d;                // put the packet to the tx fifo 
        inp_addr <= inp_addr + 1;           // increment the current pos
                                            // check the socket is matching
        if (inp_addr == 0x10)               // check the ecpri write flag is set 
        begin
            if (inp_d == 0x10) begin        // check the write flag
                send_write_resp <= 1;
            end
            if (inp_d == 0x00) begin        // check the read flag
                send_read_resp <= 1;
            end
        end
    end
end

// copy to the remote memory
always @(posedge inp_clk)
begin
if (send_write_resp) 
begin
    // get the length of the payload 
    if (inp_addr == 0x12)
    begin
        payload_len  <= inp_d;
    end

    // get the dst_address memory address 
    if (inp_addr == 0x13)
    begin
        dst_addr <= inp_d;
        tx_payload_len <= payload_len;
    end

    // copy the payload 
    if ( payload_len > 0)
    begin
        dst_addr <= inp_d;
        payload_len <= payload_len - 1;
        dst_addr <= dst_addr + 1;
    end
end

endmodule //ecpri_rx

// ram will be better option between the rx and tx module , since the 
// mac, ip & port of the src and address address has to be swapped 


/* get the data from the ram/fifo 
*/
module epcri_tx ( to_switch, data_to_mem, send_write_resp, sen_read_resp,
                    inp_clk, rx_buff, tx_payload_len, reset);

input wire reset;
input wire[7:0] rx_buff;
input wire inp_clk;
input wire out_clk;
input wire send_write_resp;
input wire read_write_resp;
output reg[7:0] to_switch;

reg [7:0] inp_addr;
integer payload_len;
integer pkt_hdr_len;

always @(posedge reset)
begin
    inp_addr <= 0;
    payload_len <= 0;
    pkt_hdr_len <= 35; //2 ip, 2 mac, 2 port, 1 vlan id, 1 ipv4 header 
end

always @(posedge clk) 
begin 
    if (send_write_resp)

    //add the mac header 
    //
    // add the ether type  
    // 
    // add the ip header 
    //
    // add the ecpri header 
    //
    // add the packet payload 
end

endmodule
